/********************************************************************
 * Model of RAM Memory - Verilog Training Course.
 *********************************************************************/

`timescale 1ns / 1ns

module mem(data,addr,read,write);
  inout [7:0] data;
  input [4:0] addr;
  input       read, write;



endmodule
