`define dly_and 1
`define dly_or 2
module mux (out,a,b,sel);





endmodule
