module rca16(sum, c_out, a, b, c_in);










endmodule
